--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:10:39 02/22/2021
-- Design Name:   
-- Module Name:   H:/Projet_Scoring/equ45min_tb.vhd
-- Project Name:  SCORING
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: equ45min
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY equ45min_tb IS
END equ45min_tb;
 
ARCHITECTURE behavior OF equ45min_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT equ45min
		Port (	min_dec : IN  std_logic_vector(3 downto 0);
				min_unit : IN  std_logic_vector(3 downto 0);
				equ : OUT  std_logic
			  );   
	END COMPONENT;
    

   --Inputs
   signal min_dec : std_logic_vector(3 downto 0) := (others => '0');
   signal min_unit : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal equ : std_logic := '0';
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: equ45min PORT MAP (
          min_dec => min_dec,
          min_unit => min_unit,
		  equ => equ
        );
		  
   -- Stimulus
   -- DUREE DU TEST : 5120ns
	 stim_proc : process
	 variable I : integer range 0 to 15 := 0;
	 variable J : integer range 0 to 15 := 0;
	 begin
		FOR I IN 0 TO 15 LOOP
			min_dec <= std_logic_vector(to_unsigned(I,4));
				FOR J IN 0 TO 15 LOOP
					min_unit <= std_logic_vector(to_unsigned(J,4));
					wait for 20ns;
				END LOOP;
		END LOOP;
      wait;
	 end process;  

END;
