----------------------------------------------------------------------------------
-- 
-- Engineer:       Renaud DAVIOT
-- 
-- Create Date:    2016 
--
-- File Name:      timeScoreFunc.vhd 
-- Module Name:    timeScoreFunc - Behavioral 
-- Project Name:   Chronoscore_VGA
--
-- Target Devices: XC3S200 (Spartan 3 - 200K)
-- 
-- Description: 
--
--
-- Revision 0.01 - File Created
--
----------------------------------------------------------------------------------

library IEEE;
    use IEEE.STD_LOGIC_1164.all;
    use IEEE.STD_LOGIC_ARITH.all;
    use IEEE.STD_LOGIC_UNSIGNED.all;

------------------------------------------------------------------------------
------------------------------------------------------------------------------

entity dataROM is 
    port (  address : in  std_logic_vector(6 downto 0);
            bitnbr  : in  std_logic_vector(1 downto 0);
            data    : out std_logic);
end dataROM;

------------------------------------------------------------------------------
------------------------------------------------------------------------------

architecture behavioral of dataROM is

--    type word     is array (0 to 3)  of std_logic;
--    type ROM_bit  is array (0 to 79) of word;
    type ROM_bit     is array (0 to 79, 0 to 3)  of std_logic;
--    type ROM_bit  is array (0 to 79) of word;
    constant bitchar: ROM_bit := (
        -- 0 --
        ('0','1','1','0'), -- 0 => 0000_000
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'), -- 7 => 0000_111

        -- 1 --
        ('0','0','1','0'), -- 8 => 0001_000
        ('0','1','1','0'),
        ('1','0','1','0'),
        ('0','0','1','0'),
        ('0','0','1','0'),
        ('0','0','1','0'),
        ('0','0','1','0'),
        ('1','1','1','1'), -- 15 => 0001_111

        -- 2 --
        ('0','1','1','0'), -- 16 => 0010_000
        ('1','0','0','1'),
        ('0','0','0','1'),
        ('0','0','1','0'),
        ('0','1','0','0'),
        ('1','0','0','0'),
        ('1','0','0','0'),
        ('0','1','1','1'), -- 23 => 0010_111

        -- 3 --
        ('0','1','1','0'), -- 24 => 0011_000
        ('1','0','0','1'),
        ('0','0','0','1'),
        ('0','1','1','1'),
        ('0','0','0','1'),
        ('0','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'), -- 31 => 0011_111

        -- 4 --
        ('0','0','1','0'), -- 32 => 0100_000
        ('0','1','1','0'),
        ('1','0','1','0'),
        ('1','0','1','0'),
        ('1','1','1','1'),
        ('0','0','1','0'),
        ('0','0','1','0'),
        ('1','1','1','1'), -- 39 => 0100_111

        -- 5 --
        ('0','1','1','1'), -- 40 => 0101_000
        ('1','0','0','0'),
        ('1','0','0','0'),
        ('1','1','0','0'),
        ('0','0','1','0'),
        ('0','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'), -- 47 => 0101_111

        -- 6 --
        ('0','0','1','1'), -- 48 => 0110_000
        ('0','1','0','0'),
        ('1','0','0','0'),
        ('1','0','0','0'),
        ('1','1','1','0'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'), -- 55 => 0110_111

        -- 7 --
        ('1','1','1','1'), -- 56 => 0111_000
        ('0','0','0','1'),
        ('0','0','1','0'),
        ('0','0','1','0'),
        ('0','1','0','0'),
        ('0','1','0','0'),
        ('0','1','0','0'),
        ('0','1','0','0'), -- 63 => 0111_111

        -- 8 --
        ('0','1','1','0'), -- 64 => 1000_000
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'),
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','0'), -- 71 => 1000_111

        -- 9 --
        ('0','1','1','0'), -- 72 => 1001_000
        ('1','0','0','1'),
        ('1','0','0','1'),
        ('0','1','1','1'),
        ('0','0','0','1'),
        ('0','0','0','1'),
        ('0','0','0','1'),
        ('1','1','1','0')  -- 79 => 1001_111
		  ); 

begin

		data <= bitchar(conv_integer(address), conv_integer(bitnbr));

end behavioral;